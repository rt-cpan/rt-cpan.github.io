`define error 1

module m ()
   wire w;

   assign w = `error;
endmodule // m
