module m ();
   wire [0:3] b;
   wire a = b[2];
endmodule
